module single (c, d, x);
input c, d;
output x;
assign x = c & d;

endmodule

