`timescale 1ns / 1ps


module alu_test;

	// Inputs
	reg [31:0]a;
	reg [31:0]b;
	reg [1:0]c;

	// Outputs
	wire [31:0]y;

	// Instantiate the Unit Under Test (UUT)
	alu uut (
		.a(a), 
		.b(b),
		.c(c), 
		.y(y)
	);

	initial begin
		// Initialize Inputs
		$dumpfile("alu_test.vcd");
     	$dumpvars(0,alu_test);
		
		 a = 32'b00101111000001001001000110000001;
		 b = 32'b01000000011100001100010001110001;
       		 c=00;
	 
	#40; 	a = 32'b10000000000000000000000001100010;
		b = 32'b00110011111111100011011110000011;	
	
	#40; 	a = 32'b00000000000000000000000000000010;
		b = 32'b11111111111111111111111111111111;
	 		

	 #40;  a = 32'b10101011111101001010101010101111;
		b = 32'b10000000001111111111110000000000;
	 #40;
	
	       a = 32'b00101111000001001001000110000001;
                 b = 32'b01000000011100001100010001110001;
                 c=01;

        #40;   a = 32'b10000000000000000000000001100010;
                b = 32'b00110011111111100011011110000011;

        #40;   a = 32'b00000000000000000000000000000010;
                b = 32'b11111111111111111111111111111111;


         #40;  a = 32'b10101011111101001010101010101111;
                b = 32'b10000000001111111111110000000000;
         #40;
		a = 32'b00101111000001001001000110000001;
                 b = 32'b01000000011100001100010001110001;
                 c=10;

        #40;   a = 32'b10000000000000000000000001100010;
                b = 32'b00110011111111100011011110000011;

        #40;   a = 32'b00000000000000000000000000000010;
                b = 32'b11111111111111111111111111111111;


         #40;  a = 32'b10101011111101001010101010101111;
                b = 32'b10000000001111111111110000000000;
         #40;
		a = 32'b00101111000001001001000110000001;
                 b = 32'b01000000011100001100010001110001;
                 c=11;

        #40;   a = 32'b10000000000000000000000001100010;
                b = 32'b00110011111111100011011110000011;

        #40;   a = 32'b00000000000000000000000000000010;
                b = 32'b11111111111111111111111111111111;


         #40;  a = 32'b10101011111101001010101010101111;
                b = 32'b10000000001111111111110000000000;
         #40;

	end
		initial begin 
		$monitor("a=%b b=%b y=%b c=%b\n",a,b,y, c);
		end
      
endmodule

